`define FIFO_DEPTH 12
`define FIFO_WIDTH 8
   
`include "interface.sv"
`include "seq_item.sv"
`include "sequence.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "scoreboard.sv"
`include "env.sv"
`include "rst_seq.sv"
`include "fifo_full_seq.sv"
`include "fifo_empty_seq.sv"
